module pctest();
wire myclk2;
clk clk2(myclk2);
PC pct(myclk2);
endmodule